`include "uvm_macros.svh"
`include "prj_pkg.svh"

module top();
    import uvm_pkg::*;
    import prj_pkg::*;

    initial
        run_test();
endmodule
